module ex_stage (
    input   wire                    clk,
    input   wire                    rst_n,
    //from id_ex_reg
    input   wire                    id_ex_reg_ALUctrl_i,
    

);