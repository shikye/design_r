module Flush_N_Branch(
    //from ex_ALU
    input   wire                    ex_branch_i,
    //to if_id_reg and id_ex_reg
    output  reg                     fnb_flush_o,
    //to id_pc
    output  reg                     fnb_jump_o
);


endmodule